module sccpu (clock, resetn, inst, pc, aluout, memeout);
input clock, resetn;
output [31:0] inst, pc, aluout, memeout;


endmodule